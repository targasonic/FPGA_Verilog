package filter_tb;

// including in order
`include "filter_driver.sv"
`include "filter_testcase.sv"
`include "filter_transaction.sv"
`include "filter_scoreboard.sv"
`include "filter_environment.sv"
`include "filter_interface.sv"
`include "filter_receiver.sv"
endpackage
