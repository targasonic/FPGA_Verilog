module filterFPGA ( clk, coefs, in, out );
		
	parameter 		IWIDTH 	= 16 ; 								//	input data (signal) width 
	parameter 		CWIDTH 	= 16 ; 								// tap coef data width (should be less then 32
	parameter 		TAPS 		= 3  ; 								//	number of filter taps

	localparam 		MWIDTH 	= (IWIDTH + CWIDTH); 			// multiplied width
	localparam 		RWIDTH 	= (MWIDTH + TAPS-1); 			// filter result width
	
	input  wire 			 					clk 	; 
	input  wire [IWIDTH 		- 1 : 0]		in  	;
	input  wire [TAPS * 16  - 1 : 0]		coefs	; 				// all input coefficient concatineted
	output wire [RWIDTH 		- 1 : 0]		out	; 				// output takes only top bits part of result

genvar i; 

generate 
	for( i = 0; i < TAPS; i = i + 1 )	
	begin:	tap 

		//make tap register chain 
		reg [IWIDTH - 1 : 0]	r	=	0 ; 
		
		if( i == 0 ) 
		begin 
			//	1 st tap takes signal from input 
			always @( posedge clk ) 
				r <= in ; 
		end 
		else 
		begin 
			//	tap reg takes signal from prev tap reg 
			always @( posedge clk ) 
				tap[i].r <= tap[i - 1].r ; 
		end 
		
		// get tap multiplication constant coef
		wire [CWIDTH - 1 : 0] c;
		assign c = coefs [ ( ( TAPS - 1 - i ) * 16 + CWIDTH - 1 ) : ( TAPS - 1 - i)* 16 ] ;
		
		//calculate multiplication and fix result in register
		reg [ MWIDTH - 1 : 0 ] m ;
		always @(posedge clk)
			m <= $signed( r ) * $signed( c );
			
		// makecombinatorial address
		reg [ MWIDTH - 1 + i : 0 ] a;
		if ( i == 0 )
		begin
			always @*
				tap [i].a = $signed ( tap[i].m );
		end
		else
		begin
			always @*
				tap [i].a = $signed ( tap[i].m ) + $signed ( tap[i- 1].a );
		end
		
	end
endgenerate


	
// fix calculate sum in register
reg [RWIDTH - 1 : 0] result ;
always @( posedge clk )
	result <= tap [TAPS - 1].a ;
	

assign out = result ;
	

endmodule